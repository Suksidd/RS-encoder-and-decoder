library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use ieee.std_logic_arith.all;  
use ieee.std_logic_unsigned.all; 

entity mul_g8 is
	port(
		clk : in STD_LOGIC;
		rst : in STD_LOGIC;		 
		m_d : in STD_LOGIC;
		a : in STD_LOGIC_VECTOR(7 downto 0);
		b : in STD_LOGIC_VECTOR(7 downto 0);
		res : out STD_LOGIC_VECTOR(7 downto 0)
		);
end mul_g8;


architecture mul_g8 of mul_g8 is
	
	component reed_sol_mull_div is
		port(
			clk : in STD_LOGIC;
			rst : in STD_LOGIC;
			a : in STD_LOGIC_VECTOR(7 downto 0);
			b : in STD_LOGIC_VECTOR(7 downto 0);	
			m_d : in STD_LOGIC;	-- '0' - mull, '1' - div
			tabla0 : in STD_LOGIC_VECTOR(7 downto 0);
			tablb0 : in STD_LOGIC_VECTOR(7 downto 0);
			tabl1 : in STD_LOGIC_VECTOR(7 downto 0);	 
			addra : out STD_LOGIC_VECTOR(7 downto 0);
			addrb : out STD_LOGIC_VECTOR(7 downto 0); 
			addr1 : out STD_LOGIC_VECTOR(7 downto 0); 
			error : out STD_LOGIC; 
			res : out STD_LOGIC_VECTOR(7 downto 0)
			);
	end component;
	
	type trom is array(0 to 255) of integer;
	constant rom0 : trom :=(						  ---2**
	1,  2,  4,  8,  16, 32, 64, 128,29, 58, 116,232,205,135,19, 38,
	76, 152,45, 90, 180,117,234,201,143,3,  6,  12, 24, 48, 96, 192,
	157,39, 78, 156,37, 74, 148,53, 106,212,181,119,238,193,159,35,
	70, 140,5,  10, 20, 40, 80, 160,93, 186,105,210,185,111,222,161,
	95, 190,97, 194,153,47, 94, 188,101,202,137,15, 30, 60, 120,240,
	253,231,211,187,107,214,177,127,254,225,223,163,91, 182,113,226,
	217,175,67, 134,17, 34, 68, 136,13, 26, 52, 104,208,189,103,206,
	129,31, 62, 124,248,237,199,147,59, 118,236,197,151,51, 102,204,
	133,23, 46, 92, 184,109,218,169,79, 158,33, 66, 132,21, 42, 84,
	168,77, 154,41, 82, 164,85, 170,73, 146,57, 114,228,213,183,115,
	230,209,191,99, 198,145,63, 126,252,229,215,179,123,246,241,255,
	227,219,171,75, 150,49, 98, 196,149,55, 110,220,165,87, 174,65,
	130,25, 50, 100,200,141,7,  14, 28, 56, 112,224,221,167,83, 166,
	81, 162,89, 178,121,242,249,239,195,155,43, 86, 172,69, 138,9,
	18, 36, 72, 144,61, 122,244,245,247,243,251,235,203,139,11, 22,
	44, 88, 176,125,250,233,207,131,27, 54, 108,216,173,71, 142,0
	); 
	constant rom1 : trom :=(					 --- log2
	255,0,  1,  25, 2,  50, 26, 198,3,  223,51, 238,27, 104,199,75,
	4,	100,224,14, 52, 141,239,129,28, 193,105,248,200,8, 76, 113,
	5,  138,101,47, 225,36, 15, 33, 53, 147,142,218,240,18, 130,69,
	29, 181,194,125,106,39, 249,185,201,154,9,  120,77, 228,114,166, 
	6,  191,139,98, 102,221,48, 253,226,152,37, 179,16, 145,34, 136,
	54, 208,148,206,143,150,219,189,241,210,19, 92, 131,56, 70, 64,
	30, 66, 182,163,195,72, 126,110,107,58, 40, 84, 250,133,186,61,
	202,94, 155,159,10, 21, 121,43, 78, 212,229,172,115,243,167,87,
	7,  112,192,247,140,128,99, 13, 103,74, 222,237,49, 197,254,24,
	227,165,153,119,38, 184,180,124,17, 68, 146,217,35, 32, 137,46,
	55, 63, 209,91, 149,188,207,205,144,135,151,178,220,252,190,97,
	242,86, 211,171,20, 42, 93, 158,132,60, 57, 83, 71, 109,65, 162,
	31, 45, 67, 216,183,123,164,118,196,23, 73, 236,127,12, 111,246,
	108,161,59, 82, 41, 157,85, 170,251,96, 134,177,187,204,62, 90,
	203,89, 95, 176,156,169,160,81, 11, 245,22, 235,122,117,44, 215,
	79, 174,213,233,230,231,173,232,116,214,244,234,168,80, 88, 175
	);	   	  	 
	
	
	signal a00,a01,a02 : std_logic_vector(7 downto 0) := (others => '0');
	signal d00,d01,d02 : std_logic_vector(7 downto 0) := (others => '0');
begin
	
	
	
	mull0: reed_sol_mull_div
	port map(
		clk => clk,
		rst => rst,
		a =>  a,	  
		b => b,
		m_d => m_d, -- mull, '1' - div
		tabla0 => d00,
		tablb0 => d01,
		tabl1  => d02,	 
		addra => a00,
		addrb => a01, 
		addr1 => a02,
		error => open, 
		res => res
		);	 	 	
	
	d00	<= conv_std_logic_vector (rom1(conv_integer(a00)),8);		 
	d01	<= conv_std_logic_vector (rom1(conv_integer(a01)),8);		 
	d02	<= conv_std_logic_vector (rom0(conv_integer(a02)),8);
	
	
	
	
end mul_g8;
